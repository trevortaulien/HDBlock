architecture RTL of SB1_1 is

    begin

    O_P0 <= '0';

end RTL;